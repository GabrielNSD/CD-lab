ENTITY SinalLO IS
PORT(a,b,c,d : IN BIT;
		S : OUT BIT);
END;
ARCHITECTURE bevah OF SinalLO IS 
COMPONENT PortaAnd2pinos IS 
PORT(en1, en2 : IN BIT;
		s0 : OUT BIT
);
END COMPONENT;
COMPONENT PortaAnd3pinos IS 
PORT(en1, en2, en3 : IN BIT;
		s0 : OUT BIT
);
END COMPONENT;
COMPONENT PortaAnd4pinos IS 
PORT(en1, en2, en3,en4 : IN BIT;
		s0 : OUT BIT
);
END COMPONENT;
COMPONENT PortaOr6pinos IS 
PORT(en1, en2, en3, en4, en5, en6  : IN BIT;
		sOr : OUT BIT
);
END COMPONENT;
SIGNAL S1: BIT;
SIGNAL S2: BIT;
SIGNAL S3: BIT;
SIGNAL S4: BIT;
SIGNAL S5: BIT;
SIGNAL S6: BIT;
BEGIN 
u1 : PortaAnd2pinos PORT MAP(en1 => not(a), en2 => not(b), s0 => S1);
u2 : PortaAnd3pinos PORT MAP(en1 => a, en2 => c, en3 => d , s0 => S2);
u3 : PortaAnd3pinos PORT MAP(en1 => not(a), en2 => b, en3 => c , s0 => S3);
u4 : PortaAnd4pinos PORT MAP(en1 => a, en2 => not(b), en3 => c , en4 => not(d), s0 => S4); 
u5 : PortaAnd4pinos PORT MAP(en1 => a, en2 => not(b), en3 => not(c) , en4 => d, s0 => S5);
u6 : PortaAnd4pinos PORT MAP(en1 => not(a), en2 => b, en3 => not(c) , en4 => d, s0 => S6);
usaida : portaOr6pinos PORT MAP(en1 => S1, en2 => S2,en3 => S3,en4 => S4,en5 => S5,en6 => S6,sOr => S);
END;
