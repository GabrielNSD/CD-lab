ENTITY Mux2x1 IS
PORT(A,B,S : IN BIT;
		X: OUT BIT);
END Mux2x1;

ARCHITECTURE Behave OF Mux2x1 IS
	SIGNAL AND1: BIT; --Recebe o sinal da primeira porta AND
	SIGNAL AND2: BIT; -- Recebe o sinal da segunda porta AND
	
	COMPONENT PortaAND IS
		PORT(AND_IN_A, AND_IN_B: IN BIT;
				AND_OUT: OUT BIT);
	END COMPONENT;
	
	COMPONENT PortaOR IS
		PORT(OR_IN_A,OR_IN_B : IN BIT;
			OR_OUT: OUT BIT);
	END COMPONENT;

BEGIN
u1: PortaAND PORT MAP(AND_IN_A=>A, AND_IN_B=>NOT S,AND_OUT=>AND1);
u2: PortaAND PORT MAP(AND_IN_A=>B, AND_IN_B=>S,AND_OUT=>AND2);
u3: PortaOR PORT MAP(OR_IN_A=>AND1,OR_IN_B=>AND2,OR_OUT=>X);
END;