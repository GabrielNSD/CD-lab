ENTITY PortaAND IS
	PORT(AND_IN_A,AND_IN_B : IN BIT;
			AND_OUT: OUT BIT);
END PortaAND;

ARCHITECTURE Behave OF PortaAND IS
BEGIN
	AND_OUT <= AND_IN_A AND AND_IN_B;
END Behave;